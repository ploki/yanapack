* SURROUND based on Fostex FF165WK and SEAS 27TFFC

.include circuits/driver.cir
.include circuits/closed_cab.cir

.subckt low_pass in out com
* filter *
Llp1 in     0  0.8m .22
Llp2  0     1  0.5m .21
Llp3  1   out  0.5m .21
Clp1  out com  12u
Clp2  out com  3.3u
* imp comp *
Cnw  out 2 1.2u
Rnw  2 com 6.8
.ends

.subckt high_pass in out com
Ratt1 in 1 5.6
Ratt2 in 1 10
Chp1 in 1 2.7u
Chp2 1 out 4.7u
Lhp out com .3m .13
*Cnt out 1 2.2u
*Rnt 1 com 4.7
.ends

* amp *
Eg 1 0 2.83

** midbass **
Xlow_pass 1 2 0 low_pass
* Fostex FF165WK *
Xmidbass 2 0 aGND 3 driver param: { .056m TO Le 6.5 TO Re 7.227 TO Bl \
			            0.7123 TO Rms 1.068m TO Cms 9.5m TO Mms \
			            132cm² TO Sd }

XBox  3 aGND closed_cab param: { 9L TO Vb 50 TO Qb 7 TO Ql \
                                 .056m TO Le 6.5 TO Re 7.227 TO Bl \
				 0.7123 TO Rms 1.068m TO Cms 9.5m TO Mms \
				 132cm² TO Sd }
*Set Vb to 15.83 to use the port
*Port  8 aGND 6.7cm 19.63cm² kKr


** tweeter **
Xhigh_pass 1 4 0 high_pass
* SEAS 27TFFC
Xtweeter 4 0 aGND aGND driver param: { .05m TO Le 4.8 TO Re 3.5 TO Bl \
                                      2 TO Rms .23m TO Cms .25m TO Mms \
	                              7.6cm² TO Sd }


* set logscale x
* set mxtics
* set mytics
* set style line 12 lc rgb '#ddccdd' lt 1 lw 1.5
* set style line 13 lc rgb '#ddccdd' lt 1 lw 0.5
* set grid xtics mxtics ytics mytics back ls 12, ls 13
* plot [16:40000] [40:100] 'plop.txt' using 1:2 title 'sum' with lines, 'plop.txt' using 1:3 title 'woofer' with lines, 'plop.txt' using 1:4 title 'tweeter' with lines

!general properties
. 132cm² TO woofer_Sd  IZfront:Xmidbass TO woofer_volume_velocity
. 7.6cm² TO tweeter_Sd IZfront:Xtweeter TO tweeter_volume_velocity
. 14.5cm TO distance_between_drivers
. 1 TO distance

!! frequency response /1m
.include circuits/frequency_response_2way.fth

!! horizontal directivity
*.include circuits/horizontal_directivity_2way.fth

!! vertical directivity
*. -5° TO vertical_angle
*.include circuits/vertical_directivity_2way.fth

! cone disp in mm
*.include circuits/cone_displacement_2way.fth

!phase
*.include circuits/phase_2way.fth

! phase delay in ms
*.include circuits/phase_delay_2way.fth

! ** group delay **
*. >>> F IZfront:Xtweeter IZfront:Xmidbass <<<
*.     TO _woofer_volume_velocity
*.     TO _tweeter_volume_velocity
*.     TO _F
*.include circuits/group_delay_2way.fth

! power dissipation in resistors
*. F .
*. IRbsc v1 v2 - * REAL ABS .
*. IRnw v4 v0 - *  REAL ABS .
*. IRatt v1 v10 - * REAL ABS .

!! power dissipation in driver's R
*. F .
*! active power
*. IEg v1 v0 - * REAL ABS .
*! reactive power
*. IEg v1 v0 - * IMAG ABS .
*! power dissipated in midbass
*. IRe:Xmidbass v0:Xmidbass v1:Xmidbass - * REAL ABS .
*! power dissipated in tweeter
*. IRe:Xtweeter v0:Xtweeter v1:Xtweeter - * REAL ABS .
*! power dissipated in the midbass suspension
**. IRrms:Xff165wk v2:Xff165wk v3:Xff165wk - * REAL ABS .
*! power dissipated in the tweeter suspension
**. IRrms:X27tffc v2:X27tffc v3:X27tffc - * REAL ABS .

! total impedance
*. F .
*. v1 v0 - IEg / DUP ABS . ARG DEG .
