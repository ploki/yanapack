* SURROUND based on Fostex FF165WK and SEAS 19TTF1

*.include driver.cir
.subckt driver in+ in- pd+ pd-
******************************
* drop: V, flow: A
Le                 in+    0   {Le}
Re                   0    1   {Re}
Glmotor              1  in-   {1 Bl /}
Rmotor_linkage     in-    g   1T
Grmotor              2    g   {1 Bl /}
* drop: N, flow: m/s
Rrms                 2    3   {Rms}
Lmms                 3    4   {Mms}
Ccms                 4    5   {Cms}
Tldiaphragm          5    g   {Sd}
Rdiaphragm_linkage   g  pd-   1T
Trdiaphragm        pd+  pd-   1
* drop: Pa, flow: m³/s
.ends

* amp *
Eg 1 0 2.83

** midbass **

* bsc *
Lbsc 1 2 0.8m .22
Rbsc 1 2 3.3

* low pass *
Llp  2 3 .6m .21
Clp  3 0 5.6u

* imp comp *
Cnw  3 4 1.2u
Rnw  4 0 6.8

* driver *
Xff165wk 3 0 7 5 driver param: { .056m TO Le 6.5 TO Re 7.227 TO Bl \
			         0.7123 TO Rms 1.068m TO Cms 9.5m TO Mms \
			         132cm² TO Sd }

ZrW1  7 8 132cm² ai
Box   8 9 9L
ZrWr  9 5 132cm² ai

** tweeter **

Ratt 1 10 5.6
Chp 10 11 3.3u
Lhp 11 0 .15m .09

*Cnt 11 12 2.2u
*Rnt 12 0 4.7

X27tffc 11 0 15 13 driver param: { .05m TO Le 4.8 TO Re 3.5 TO Bl \
                                   2 TO Rms .23m TO Cms .25m TO Mms \
	                           7.6cm² TO Sd }
ZrT1  15 16 7.6cm² ai
ZrT2  16 13 7.6cm² ai


* set logscale x
* set mxtics
* set mytics
* set style line 12 lc rgb '#ddccdd' lt 1 lw 1.5
* set style line 13 lc rgb '#ddccdd' lt 1 lw 0.5
* set grid xtics mxtics ytics mytics back ls 12, ls 13
* plot [16:40000] [40:100] 'plop.txt' using 1:2 title 'sum' with lines, 'plop.txt' using 1:3 title 'woofer' with lines, 'plop.txt' using 1:4 title 'tweeter' with lines

! frequency response /1m
. F .
. 132cm² 1 0° DIRIMP IZrW1 * 7.6cm² 1 0° DIRIMP IZrT1 * - DBSPL .
. 132cm² 1 0° DIRIMP IZrW1 * DBSPL .
. 7.6cm² 1 0° DIRIMP IZrT1 * DBSPL .

*. F . 
*. 132cm² 1 0° DIRIMP IZrW1 *
*. 7.6cm² 1 0° DIRIMP IZrT1 * - DBSPL .
*. 132cm² 1 30° DIRIMP IZrW1 *
*. 7.6cm² 1 30° DIRIMP IZrT1 * - DBSPL .
*. 132cm² 1 60° DIRIMP IZrW1 *
*. 7.6cm² 1 60° DIRIMP IZrT1 * - DBSPL .


! cone disp
*. F .
*. IZrW1 ABS 2 SQRT * 2 PI * F * 132cm² * / 1000 * .


!phase
*. F .
*. IZrW1 ARG .
*. IZrT1 ARG .

! power dissipation in resistors
*. F .
*. IRbsc v1 v2 - * REAL ABS .
*. IRnw v4 v0 - *  REAL ABS .

! total impedance
*. F .
*. v1 v0 - IEg / DUP ABS . ARG DEG .

! phase delay
*. F DUP .
*. 1 SWAP / 1000 * DUP NEG . .
*. 
*. IZrW1 ARG PDELAY 1000 * .
*. IZrT1 ARG PDELAY 1000 * .
*. IZrW1 ARG .

! ** group delay **
*. >>> F <<< F - 2 PI * * 1000 /
*. DUP
*! freq
*. F DUP .
*! -1 cycle and 1 cycle
*. 1 SWAP / 1000 * DUP NEG . .
*! group delay of the midbass driver
*. >>> IZrW1 ARG <<< IZrW1 ARG ANGLE SWAP / NEG .
*! group delay of the HF driver
*. >>> IZrT1 ARG <<< IZrT1 ARG ANGLE SWAP / NEG .
*! phase of the midbass driver
*. IZrW1 ARG .
